module mux16_1 (
    input logic [3:0] sel,
    input logic [15:0] d,
    output logic q,
);
// first stage of four
// generate four 

endmodule