module DFF_enable (
    output logic q;
    input logic d, reset, clk, enable;
);

endmodule