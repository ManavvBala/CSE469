module CPU (
    input logic clock,
    input logic reset
);
    

endmodule